library verilog;
use verilog.vl_types.all;
entity trans3to8_vlg_vec_tst is
end trans3to8_vlg_vec_tst;
